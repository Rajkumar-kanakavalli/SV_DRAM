/* package ram_pkg;

   int number_of_transactions=1;
   
   `include "transaction.sv"
   `include "generator.sv"
   `include "write_driver.sv"
   `include "read_driver.sv"
   `include "write_monitor.sv"
   `include "read_monitor.sv"
   `include "reference_model.sv"
   `include "scoreboard.sv"
   `include "environment.sv"
   
   endpackage */